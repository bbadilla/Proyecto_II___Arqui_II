module Add_pc(input logic [17:0] a, input logic [17:0] b,
				output logic [17:0] c);
	
	assign c = a + b;

endmodule
