module acumulator(input logic clk, we, input logic [15:0] ram[255:0], output logic [127:0] out_ac);
	
	logic [15:0] mem[255:0];
	logic [15:0] adder_out [254:0];
	Add_param #(16) add_ac(ram[0], ram[1], adder_out[0]);

	
	genvar i;
	generate
		for(i = 1; i < 255; i++)
		begin:ac
			Add_param #(16) add_ac(adder_out[i - 1], ram[i + 1], adder_out[i]);
		end
	endgenerate
	
	generate
		 for(i = 0; i < 256; i++)
		 begin: test
			  initial
			  begin
					mem[i][15:0] = 16'b0;
			  end
		 end
	endgenerate
	
	always_ff @(posedge clk)
    if (we)
		begin
			mem[0] <= ram[0];  
			mem[1] <= adder_out[0];
			mem[2] <= adder_out[1];
			mem[3] <= adder_out[2];
			mem[4] <= adder_out[3];
			mem[5] <= adder_out[4];
			mem[6] <= adder_out[5];
			mem[7] <= adder_out[6];
			mem[8] <= adder_out[7];
			mem[9] <= adder_out[8];
			mem[10] <= adder_out[9];
			mem[11] <= adder_out[10];
			mem[12] <= adder_out[11];
			mem[13] <= adder_out[12];
			mem[14] <= adder_out[13];
			mem[15] <= adder_out[14];
			mem[16] <= adder_out[15];
			mem[17] <= adder_out[16];
			mem[18] <= adder_out[17];
			mem[19] <= adder_out[18];
			mem[20] <= adder_out[19];
			mem[21] <= adder_out[20];
			mem[22] <= adder_out[21];
			mem[23] <= adder_out[22];
			mem[24] <= adder_out[23];
			mem[25] <= adder_out[24];
			mem[26] <= adder_out[25];
			mem[27] <= adder_out[26];
			mem[28] <= adder_out[27];
			mem[29] <= adder_out[28];
			mem[30] <= adder_out[29];
			mem[31] <= adder_out[30];
			mem[32] <= adder_out[31];
			mem[33] <= adder_out[32];
			mem[34] <= adder_out[33];
			mem[35] <= adder_out[34];
			mem[36] <= adder_out[35];
			mem[37] <= adder_out[36];
			mem[38] <= adder_out[37];
			mem[39] <= adder_out[38];
			mem[40] <= adder_out[39];
			mem[41] <= adder_out[40];
			mem[42] <= adder_out[41];
			mem[43] <= adder_out[42];
			mem[44] <= adder_out[43];
			mem[45] <= adder_out[44];
			mem[46] <= adder_out[45];
			mem[47] <= adder_out[46];
			mem[48] <= adder_out[47];
			mem[49] <= adder_out[48];
			mem[50] <= adder_out[49];
			mem[51] <= adder_out[50];
			mem[52] <= adder_out[51];
			mem[53] <= adder_out[52];
			mem[54] <= adder_out[53];
			mem[55] <= adder_out[54];
			mem[56] <= adder_out[55];
			mem[57] <= adder_out[56];
			mem[58] <= adder_out[57];
			mem[59] <= adder_out[58];
			mem[60] <= adder_out[59];
			mem[61] <= adder_out[60];
			mem[62] <= adder_out[61];
			mem[63] <= adder_out[62];
			mem[64] <= adder_out[63];
			mem[65] <= adder_out[64];
			mem[66] <= adder_out[65];
			mem[67] <= adder_out[66];
			mem[68] <= adder_out[67];
			mem[69] <= adder_out[68];
			mem[70] <= adder_out[69];
			mem[71] <= adder_out[70];
			mem[72] <= adder_out[71];
			mem[73] <= adder_out[72];
			mem[74] <= adder_out[73];
			mem[75] <= adder_out[74];
			mem[76] <= adder_out[75];
			mem[77] <= adder_out[76];
			mem[78] <= adder_out[77];
			mem[79] <= adder_out[78];
			mem[80] <= adder_out[79];
			mem[81] <= adder_out[80];
			mem[82] <= adder_out[81];
			mem[83] <= adder_out[82];
			mem[84] <= adder_out[83];
			mem[85] <= adder_out[84];
			mem[86] <= adder_out[85];
			mem[87] <= adder_out[86];
			mem[88] <= adder_out[87];
			mem[89] <= adder_out[88];
			mem[90] <= adder_out[89];
			mem[91] <= adder_out[90];
			mem[92] <= adder_out[91];
			mem[93] <= adder_out[92];
			mem[94] <= adder_out[93];
			mem[95] <= adder_out[94];
			mem[96] <= adder_out[95];
			mem[97] <= adder_out[96];
			mem[98] <= adder_out[97];
			mem[99] <= adder_out[98];
			mem[100] <= adder_out[99];
			mem[101] <= adder_out[100];
			mem[102] <= adder_out[101];
			mem[103] <= adder_out[102];
			mem[104] <= adder_out[103];
			mem[105] <= adder_out[104];
			mem[106] <= adder_out[105];
			mem[107] <= adder_out[106];
			mem[108] <= adder_out[107];
			mem[109] <= adder_out[108];
			mem[110] <= adder_out[109];
			mem[111] <= adder_out[110];
			mem[112] <= adder_out[111];
			mem[113] <= adder_out[112];
			mem[114] <= adder_out[113];
			mem[115] <= adder_out[114];
			mem[116] <= adder_out[115];
			mem[117] <= adder_out[116];
			mem[118] <= adder_out[117];
			mem[119] <= adder_out[118];
			mem[120] <= adder_out[119];
			mem[121] <= adder_out[120];
			mem[122] <= adder_out[121];
			mem[123] <= adder_out[122];
			mem[124] <= adder_out[123];
			mem[125] <= adder_out[124];
			mem[126] <= adder_out[125];
			mem[127] <= adder_out[126];
			mem[128] <= adder_out[127];
			mem[129] <= adder_out[128];
			mem[130] <= adder_out[129];
			mem[131] <= adder_out[130];
			mem[132] <= adder_out[131];
			mem[133] <= adder_out[132];
			mem[134] <= adder_out[133];
			mem[135] <= adder_out[134];
			mem[136] <= adder_out[135];
			mem[137] <= adder_out[136];
			mem[138] <= adder_out[137];
			mem[139] <= adder_out[138];
			mem[140] <= adder_out[139];
			mem[141] <= adder_out[140];
			mem[142] <= adder_out[141];
			mem[143] <= adder_out[142];
			mem[144] <= adder_out[143];
			mem[145] <= adder_out[144];
			mem[146] <= adder_out[145];
			mem[147] <= adder_out[146];
			mem[148] <= adder_out[147];
			mem[149] <= adder_out[148];
			mem[150] <= adder_out[149];
			mem[151] <= adder_out[150];
			mem[152] <= adder_out[151];
			mem[153] <= adder_out[152];
			mem[154] <= adder_out[153];
			mem[155] <= adder_out[154];
			mem[156] <= adder_out[155];
			mem[157] <= adder_out[156];
			mem[158] <= adder_out[157];
			mem[159] <= adder_out[158];
			mem[160] <= adder_out[159];
			mem[161] <= adder_out[160];
			mem[162] <= adder_out[161];
			mem[163] <= adder_out[162];
			mem[164] <= adder_out[163];
			mem[165] <= adder_out[164];
			mem[166] <= adder_out[165];
			mem[167] <= adder_out[166];
			mem[168] <= adder_out[167];
			mem[169] <= adder_out[168];
			mem[170] <= adder_out[169];
			mem[171] <= adder_out[170];
			mem[172] <= adder_out[171];
			mem[173] <= adder_out[172];
			mem[174] <= adder_out[173];
			mem[175] <= adder_out[174];
			mem[176] <= adder_out[175];
			mem[177] <= adder_out[176];
			mem[178] <= adder_out[177];
			mem[179] <= adder_out[178];
			mem[180] <= adder_out[179];
			mem[181] <= adder_out[180];
			mem[182] <= adder_out[181];
			mem[183] <= adder_out[182];
			mem[184] <= adder_out[183];
			mem[185] <= adder_out[184];
			mem[186] <= adder_out[185];
			mem[187] <= adder_out[186];
			mem[188] <= adder_out[187];
			mem[189] <= adder_out[188];
			mem[190] <= adder_out[189];
			mem[191] <= adder_out[190];
			mem[192] <= adder_out[191];
			mem[193] <= adder_out[192];
			mem[194] <= adder_out[193];
			mem[195] <= adder_out[194];
			mem[196] <= adder_out[195];
			mem[197] <= adder_out[196];
			mem[198] <= adder_out[197];
			mem[199] <= adder_out[198];
			mem[200] <= adder_out[199];
			mem[201] <= adder_out[200];
			mem[202] <= adder_out[201];
			mem[203] <= adder_out[202];
			mem[204] <= adder_out[203];
			mem[205] <= adder_out[204];
			mem[206] <= adder_out[205];
			mem[207] <= adder_out[206];
			mem[208] <= adder_out[207];
			mem[209] <= adder_out[208];
			mem[210] <= adder_out[209];
			mem[211] <= adder_out[210];
			mem[212] <= adder_out[211];
			mem[213] <= adder_out[212];
			mem[214] <= adder_out[213];
			mem[215] <= adder_out[214];
			mem[216] <= adder_out[215];
			mem[217] <= adder_out[216];
			mem[218] <= adder_out[217];
			mem[219] <= adder_out[218];
			mem[220] <= adder_out[219];
			mem[221] <= adder_out[220];
			mem[222] <= adder_out[221];
			mem[223] <= adder_out[222];
			mem[224] <= adder_out[223];
			mem[225] <= adder_out[224];
			mem[226] <= adder_out[225];
			mem[227] <= adder_out[226];
			mem[228] <= adder_out[227];
			mem[229] <= adder_out[228];
			mem[230] <= adder_out[229];
			mem[231] <= adder_out[230];
			mem[232] <= adder_out[231];
			mem[233] <= adder_out[232];
			mem[234] <= adder_out[233];
			mem[235] <= adder_out[234];
			mem[236] <= adder_out[235];
			mem[237] <= adder_out[236];
			mem[238] <= adder_out[237];
			mem[239] <= adder_out[238];
			mem[240] <= adder_out[239];
			mem[241] <= adder_out[240];
			mem[242] <= adder_out[241];
			mem[243] <= adder_out[242];
			mem[244] <= adder_out[243];
			mem[245] <= adder_out[244];
			mem[246] <= adder_out[245];
			mem[247] <= adder_out[246];
			mem[248] <= adder_out[247];
			mem[249] <= adder_out[248];
			mem[250] <= adder_out[249];
			mem[251] <= adder_out[250];
			mem[252] <= adder_out[251];
			mem[253] <= adder_out[252];
			mem[254] <= adder_out[253];
			mem[255] <= adder_out[254];

		end	
endmodule 