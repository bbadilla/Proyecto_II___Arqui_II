module Add (input logic [127:0] a, input logic [127:0] b,
				output logic [127:0] c);
	
	assign c = a + b;
		
endmodule
